module SingleCycle(
);

endmodule
