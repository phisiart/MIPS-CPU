module REG(
    input wire RegRd,
    input wire RegWr,
    input wire[1:0] RegDst,
    input wire[4:0] Rs,
    input wire[4:0] Rt,
    input wire[4:0] Rd,
);

    

    

endmodule
