`timescale 1ns / 1ps

// ZHENGRONG WANG
// Created 11/07/2014
// Last Modified 11/07/2014

module MEM_REG_REG(
    );


endmodule
